----------------------------------------------------------------------------------
-- CMS Muon Endcap
-- GEM Collaboration
-- Optohybrid v3 Firmware -- TDC
-- 2018/07/11 -- Initial
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.types_pkg.all;
use work.param_pkg.all;
use work.ipbus_pkg.all;
use work.registers.all;

entity oh_tdc is
port(

    -- Clocks
    clk_1x_i : in std_logic;
    clk_8x_i : in std_logic;

    -- Config
    reset_i       : in std_logic;

    -- Inputs
    trigger_i   : in std_logic;
    sbits_i     : in std_logic_vector(23 downto 0);

    -- ipbus

    ipb_mosi_i : in  ipb_wbus;
    ipb_miso_o : out ipb_rbus;

    ipb_reset_i : in std_logic;
    ipb_clk_i : in std_logic

);
end oh_tdc;


architecture Behavioral of oh_tdc is

    signal reset : std_logic;
    signal reset_local : std_logic;
    signal resetting : std_logic;

    signal calibrate : std_logic;
    signal calibrating : std_logic;
    signal window_mask : std_logic_vector (255 downto 0);
    signal vfat_mask : std_logic_vector (23 downto 0);
    signal fifo_rden : std_logic_vector (23 downto 0);
    signal fifo_dout : std32_array_t (23 downto 0);
    signal fifo_valid : std_logic_vector (23 downto 0);
    signal callut_addr : std_logic_vector(8 downto 0);
    signal callut_data : std_logic_vector(11 downto 0);

    signal callut_addr_pulse, callut_addr_progress, callut_addr_done : std_logic;

    ------ Register signals begin (this section is generated by <optohybrid_top>/tools/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_TDC_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------

begin

    process (clk_1x_i) begin
        if (rising_edge(clk_1x_i)) then
            reset <= reset_local or reset_i;
        end if;
    end process;

    tdc_inst : entity work.tdc
    port map (
        clk_1x_i => clk_1x_i,
        clk_8x_i => clk_8x_i,

        -- Config
        reset_i       => reset,
        resetting_o   => resetting,

        calibrate_i   => calibrate,
        calibrating_o => calibrating,

        window_mask_i => window_mask,
        vfat_mask_i   => vfat_mask,

        -- Inputs
        trigger_i  => trigger_i,
        sbits_i    => sbits_i,

        -- FIFOs
        fifo_rden      => fifo_rden,
        fifo_dout      => fifo_dout,
        fifo_valid     => fifo_valid,
        fifo_underflow => open,

        -- Calibration LUT
        callut_addr_i => callut_addr,
        callut_data_o => callut_data

    );

    -- Delay the address write of two clock cycles to be sure to read the correct data on the next read
    process(clk_1x_i) begin
        if (rising_edge(clk_1x_i)) then
            callut_addr_done     <= callut_addr_progress;
            callut_addr_progress <= callut_addr_pulse;
        end if;
    end process;

    --===============================================================================================
    -- (this section is generated by <optohybrid_top>/tools/generate_registers.py -- do not edit)
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_TDC_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_TDC_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_TDC_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clk_1x_i,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"0";
    regs_addresses(1)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"1";
    regs_addresses(2)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"2";
    regs_addresses(3)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"3";
    regs_addresses(4)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"4";
    regs_addresses(5)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"5";
    regs_addresses(6)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"6";
    regs_addresses(7)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"7";
    regs_addresses(8)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"8";
    regs_addresses(9)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"9";
    regs_addresses(10)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"a";
    regs_addresses(11)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"b";
    regs_addresses(12)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"c";
    regs_addresses(13)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"d";
    regs_addresses(14)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"0";
    regs_addresses(15)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"1";
    regs_addresses(16)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"2";
    regs_addresses(17)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"3";
    regs_addresses(18)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"4";
    regs_addresses(19)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"5";
    regs_addresses(20)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"6";
    regs_addresses(21)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"7";
    regs_addresses(22)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"8";
    regs_addresses(23)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"9";
    regs_addresses(24)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"a";
    regs_addresses(25)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"b";
    regs_addresses(26)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"c";
    regs_addresses(27)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"d";
    regs_addresses(28)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"e";
    regs_addresses(29)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"f";
    regs_addresses(30)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "11" & x"0";
    regs_addresses(31)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "11" & x"1";
    regs_addresses(32)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "11" & x"2";
    regs_addresses(33)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "11" & x"3";
    regs_addresses(34)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "11" & x"4";
    regs_addresses(35)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "11" & x"5";
    regs_addresses(36)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "11" & x"6";
    regs_addresses(37)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "11" & x"7";

    -- Connect read signals
    regs_read_arr(1)(REG_TDC_CTRL_RESETTING_BIT) <= resetting;
    regs_read_arr(3)(REG_TDC_CTRL_CALIBRATING_BIT) <= calibrating;
    regs_read_arr(4)(REG_TDC_CTRL_CALLUT_DATA_MSB downto REG_TDC_CTRL_CALLUT_DATA_LSB) <= callut_data;
    regs_read_arr(4)(REG_TDC_CTRL_CALLUT_ADDR_MSB downto REG_TDC_CTRL_CALLUT_ADDR_LSB) <= callut_addr;
    regs_read_arr(5)(REG_TDC_CTRL_VFAT_MASK_MSB downto REG_TDC_CTRL_VFAT_MASK_LSB) <= vfat_mask;
    regs_read_arr(6)(REG_TDC_CTRL_WINDOW_MASK_0_MSB downto REG_TDC_CTRL_WINDOW_MASK_0_LSB) <= window_mask(31 downto 0);
    regs_read_arr(7)(REG_TDC_CTRL_WINDOW_MASK_1_MSB downto REG_TDC_CTRL_WINDOW_MASK_1_LSB) <= window_mask(63 downto 32);
    regs_read_arr(8)(REG_TDC_CTRL_WINDOW_MASK_2_MSB downto REG_TDC_CTRL_WINDOW_MASK_2_LSB) <= window_mask(95 downto 64);
    regs_read_arr(9)(REG_TDC_CTRL_WINDOW_MASK_3_MSB downto REG_TDC_CTRL_WINDOW_MASK_3_LSB) <= window_mask(127 downto 96);
    regs_read_arr(10)(REG_TDC_CTRL_WINDOW_MASK_4_MSB downto REG_TDC_CTRL_WINDOW_MASK_4_LSB) <= window_mask(159 downto 128);
    regs_read_arr(11)(REG_TDC_CTRL_WINDOW_MASK_5_MSB downto REG_TDC_CTRL_WINDOW_MASK_5_LSB) <= window_mask(191 downto 160);
    regs_read_arr(12)(REG_TDC_CTRL_WINDOW_MASK_6_MSB downto REG_TDC_CTRL_WINDOW_MASK_6_LSB) <= window_mask(223 downto 192);
    regs_read_arr(13)(REG_TDC_CTRL_WINDOW_MASK_7_MSB downto REG_TDC_CTRL_WINDOW_MASK_7_LSB) <= window_mask(255 downto 224);
    regs_read_arr(14)(REG_TDC_FIFOS_VFAT0_MSB downto REG_TDC_FIFOS_VFAT0_LSB) <= fifo_dout(0);
    regs_read_arr(15)(REG_TDC_FIFOS_VFAT1_MSB downto REG_TDC_FIFOS_VFAT1_LSB) <= fifo_dout(1);
    regs_read_arr(16)(REG_TDC_FIFOS_VFAT2_MSB downto REG_TDC_FIFOS_VFAT2_LSB) <= fifo_dout(2);
    regs_read_arr(17)(REG_TDC_FIFOS_VFAT3_MSB downto REG_TDC_FIFOS_VFAT3_LSB) <= fifo_dout(3);
    regs_read_arr(18)(REG_TDC_FIFOS_VFAT4_MSB downto REG_TDC_FIFOS_VFAT4_LSB) <= fifo_dout(4);
    regs_read_arr(19)(REG_TDC_FIFOS_VFAT5_MSB downto REG_TDC_FIFOS_VFAT5_LSB) <= fifo_dout(5);
    regs_read_arr(20)(REG_TDC_FIFOS_VFAT6_MSB downto REG_TDC_FIFOS_VFAT6_LSB) <= fifo_dout(6);
    regs_read_arr(21)(REG_TDC_FIFOS_VFAT7_MSB downto REG_TDC_FIFOS_VFAT7_LSB) <= fifo_dout(7);
    regs_read_arr(22)(REG_TDC_FIFOS_VFAT8_MSB downto REG_TDC_FIFOS_VFAT8_LSB) <= fifo_dout(8);
    regs_read_arr(23)(REG_TDC_FIFOS_VFAT9_MSB downto REG_TDC_FIFOS_VFAT9_LSB) <= fifo_dout(9);
    regs_read_arr(24)(REG_TDC_FIFOS_VFAT10_MSB downto REG_TDC_FIFOS_VFAT10_LSB) <= fifo_dout(10);
    regs_read_arr(25)(REG_TDC_FIFOS_VFAT11_MSB downto REG_TDC_FIFOS_VFAT11_LSB) <= fifo_dout(11);
    regs_read_arr(26)(REG_TDC_FIFOS_VFAT12_MSB downto REG_TDC_FIFOS_VFAT12_LSB) <= fifo_dout(12);
    regs_read_arr(27)(REG_TDC_FIFOS_VFAT13_MSB downto REG_TDC_FIFOS_VFAT13_LSB) <= fifo_dout(13);
    regs_read_arr(28)(REG_TDC_FIFOS_VFAT14_MSB downto REG_TDC_FIFOS_VFAT14_LSB) <= fifo_dout(14);
    regs_read_arr(29)(REG_TDC_FIFOS_VFAT15_MSB downto REG_TDC_FIFOS_VFAT15_LSB) <= fifo_dout(15);
    regs_read_arr(30)(REG_TDC_FIFOS_VFAT16_MSB downto REG_TDC_FIFOS_VFAT16_LSB) <= fifo_dout(16);
    regs_read_arr(31)(REG_TDC_FIFOS_VFAT17_MSB downto REG_TDC_FIFOS_VFAT17_LSB) <= fifo_dout(17);
    regs_read_arr(32)(REG_TDC_FIFOS_VFAT18_MSB downto REG_TDC_FIFOS_VFAT18_LSB) <= fifo_dout(18);
    regs_read_arr(33)(REG_TDC_FIFOS_VFAT19_MSB downto REG_TDC_FIFOS_VFAT19_LSB) <= fifo_dout(19);
    regs_read_arr(34)(REG_TDC_FIFOS_VFAT20_MSB downto REG_TDC_FIFOS_VFAT20_LSB) <= fifo_dout(20);
    regs_read_arr(35)(REG_TDC_FIFOS_VFAT21_MSB downto REG_TDC_FIFOS_VFAT21_LSB) <= fifo_dout(21);
    regs_read_arr(36)(REG_TDC_FIFOS_VFAT22_MSB downto REG_TDC_FIFOS_VFAT22_LSB) <= fifo_dout(22);
    regs_read_arr(37)(REG_TDC_FIFOS_VFAT23_MSB downto REG_TDC_FIFOS_VFAT23_LSB) <= fifo_dout(23);

    -- Connect write signals
    callut_addr <= regs_write_arr(4)(REG_TDC_CTRL_CALLUT_ADDR_MSB downto REG_TDC_CTRL_CALLUT_ADDR_LSB);
    vfat_mask <= regs_write_arr(5)(REG_TDC_CTRL_VFAT_MASK_MSB downto REG_TDC_CTRL_VFAT_MASK_LSB);
    window_mask(31 downto 0) <= regs_write_arr(6)(REG_TDC_CTRL_WINDOW_MASK_0_MSB downto REG_TDC_CTRL_WINDOW_MASK_0_LSB);
    window_mask(63 downto 32) <= regs_write_arr(7)(REG_TDC_CTRL_WINDOW_MASK_1_MSB downto REG_TDC_CTRL_WINDOW_MASK_1_LSB);
    window_mask(95 downto 64) <= regs_write_arr(8)(REG_TDC_CTRL_WINDOW_MASK_2_MSB downto REG_TDC_CTRL_WINDOW_MASK_2_LSB);
    window_mask(127 downto 96) <= regs_write_arr(9)(REG_TDC_CTRL_WINDOW_MASK_3_MSB downto REG_TDC_CTRL_WINDOW_MASK_3_LSB);
    window_mask(159 downto 128) <= regs_write_arr(10)(REG_TDC_CTRL_WINDOW_MASK_4_MSB downto REG_TDC_CTRL_WINDOW_MASK_4_LSB);
    window_mask(191 downto 160) <= regs_write_arr(11)(REG_TDC_CTRL_WINDOW_MASK_5_MSB downto REG_TDC_CTRL_WINDOW_MASK_5_LSB);
    window_mask(223 downto 192) <= regs_write_arr(12)(REG_TDC_CTRL_WINDOW_MASK_6_MSB downto REG_TDC_CTRL_WINDOW_MASK_6_LSB);
    window_mask(255 downto 224) <= regs_write_arr(13)(REG_TDC_CTRL_WINDOW_MASK_7_MSB downto REG_TDC_CTRL_WINDOW_MASK_7_LSB);

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);
    calibrate <= regs_write_pulse_arr(2);
    callut_addr_pulse <= regs_write_pulse_arr(4);

    -- Connect write done signals
    regs_write_done_arr(4) <= callut_addr_done;

    -- Connect read pulse signals
    fifo_rden(0) <= regs_read_pulse_arr(14);
    fifo_rden(1) <= regs_read_pulse_arr(15);
    fifo_rden(2) <= regs_read_pulse_arr(16);
    fifo_rden(3) <= regs_read_pulse_arr(17);
    fifo_rden(4) <= regs_read_pulse_arr(18);
    fifo_rden(5) <= regs_read_pulse_arr(19);
    fifo_rden(6) <= regs_read_pulse_arr(20);
    fifo_rden(7) <= regs_read_pulse_arr(21);
    fifo_rden(8) <= regs_read_pulse_arr(22);
    fifo_rden(9) <= regs_read_pulse_arr(23);
    fifo_rden(10) <= regs_read_pulse_arr(24);
    fifo_rden(11) <= regs_read_pulse_arr(25);
    fifo_rden(12) <= regs_read_pulse_arr(26);
    fifo_rden(13) <= regs_read_pulse_arr(27);
    fifo_rden(14) <= regs_read_pulse_arr(28);
    fifo_rden(15) <= regs_read_pulse_arr(29);
    fifo_rden(16) <= regs_read_pulse_arr(30);
    fifo_rden(17) <= regs_read_pulse_arr(31);
    fifo_rden(18) <= regs_read_pulse_arr(32);
    fifo_rden(19) <= regs_read_pulse_arr(33);
    fifo_rden(20) <= regs_read_pulse_arr(34);
    fifo_rden(21) <= regs_read_pulse_arr(35);
    fifo_rden(22) <= regs_read_pulse_arr(36);
    fifo_rden(23) <= regs_read_pulse_arr(37);

    -- Connect counter instances

    -- Connect rate instances

    -- Connect read ready signals
    regs_read_ready_arr(14) <= fifo_valid(0);
    regs_read_ready_arr(15) <= fifo_valid(1);
    regs_read_ready_arr(16) <= fifo_valid(2);
    regs_read_ready_arr(17) <= fifo_valid(3);
    regs_read_ready_arr(18) <= fifo_valid(4);
    regs_read_ready_arr(19) <= fifo_valid(5);
    regs_read_ready_arr(20) <= fifo_valid(6);
    regs_read_ready_arr(21) <= fifo_valid(7);
    regs_read_ready_arr(22) <= fifo_valid(8);
    regs_read_ready_arr(23) <= fifo_valid(9);
    regs_read_ready_arr(24) <= fifo_valid(10);
    regs_read_ready_arr(25) <= fifo_valid(11);
    regs_read_ready_arr(26) <= fifo_valid(12);
    regs_read_ready_arr(27) <= fifo_valid(13);
    regs_read_ready_arr(28) <= fifo_valid(14);
    regs_read_ready_arr(29) <= fifo_valid(15);
    regs_read_ready_arr(30) <= fifo_valid(16);
    regs_read_ready_arr(31) <= fifo_valid(17);
    regs_read_ready_arr(32) <= fifo_valid(18);
    regs_read_ready_arr(33) <= fifo_valid(19);
    regs_read_ready_arr(34) <= fifo_valid(20);
    regs_read_ready_arr(35) <= fifo_valid(21);
    regs_read_ready_arr(36) <= fifo_valid(22);
    regs_read_ready_arr(37) <= fifo_valid(23);

    -- Defaults
    regs_defaults(4)(REG_TDC_CTRL_CALLUT_ADDR_MSB downto REG_TDC_CTRL_CALLUT_ADDR_LSB) <= REG_TDC_CTRL_CALLUT_ADDR_DEFAULT;
    regs_defaults(5)(REG_TDC_CTRL_VFAT_MASK_MSB downto REG_TDC_CTRL_VFAT_MASK_LSB) <= REG_TDC_CTRL_VFAT_MASK_DEFAULT;
    regs_defaults(6)(REG_TDC_CTRL_WINDOW_MASK_0_MSB downto REG_TDC_CTRL_WINDOW_MASK_0_LSB) <= REG_TDC_CTRL_WINDOW_MASK_0_DEFAULT;
    regs_defaults(7)(REG_TDC_CTRL_WINDOW_MASK_1_MSB downto REG_TDC_CTRL_WINDOW_MASK_1_LSB) <= REG_TDC_CTRL_WINDOW_MASK_1_DEFAULT;
    regs_defaults(8)(REG_TDC_CTRL_WINDOW_MASK_2_MSB downto REG_TDC_CTRL_WINDOW_MASK_2_LSB) <= REG_TDC_CTRL_WINDOW_MASK_2_DEFAULT;
    regs_defaults(9)(REG_TDC_CTRL_WINDOW_MASK_3_MSB downto REG_TDC_CTRL_WINDOW_MASK_3_LSB) <= REG_TDC_CTRL_WINDOW_MASK_3_DEFAULT;
    regs_defaults(10)(REG_TDC_CTRL_WINDOW_MASK_4_MSB downto REG_TDC_CTRL_WINDOW_MASK_4_LSB) <= REG_TDC_CTRL_WINDOW_MASK_4_DEFAULT;
    regs_defaults(11)(REG_TDC_CTRL_WINDOW_MASK_5_MSB downto REG_TDC_CTRL_WINDOW_MASK_5_LSB) <= REG_TDC_CTRL_WINDOW_MASK_5_DEFAULT;
    regs_defaults(12)(REG_TDC_CTRL_WINDOW_MASK_6_MSB downto REG_TDC_CTRL_WINDOW_MASK_6_LSB) <= REG_TDC_CTRL_WINDOW_MASK_6_DEFAULT;
    regs_defaults(13)(REG_TDC_CTRL_WINDOW_MASK_7_MSB downto REG_TDC_CTRL_WINDOW_MASK_7_LSB) <= REG_TDC_CTRL_WINDOW_MASK_7_DEFAULT;

    -- Define writable regs
    regs_writable_arr(4) <= '1';
    regs_writable_arr(5) <= '1';
    regs_writable_arr(6) <= '1';
    regs_writable_arr(7) <= '1';
    regs_writable_arr(8) <= '1';
    regs_writable_arr(9) <= '1';
    regs_writable_arr(10) <= '1';
    regs_writable_arr(11) <= '1';
    regs_writable_arr(12) <= '1';
    regs_writable_arr(13) <= '1';

    --==== Registers end ============================================================================

end Behavioral;
